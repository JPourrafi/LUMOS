`include "Defines.vh"

module Fixed_Point_Unit 
#(
    parameter WIDTH = 32,
    parameter FBITS = 10
)
(
    input wire clk,
    input wire reset,
    
    input wire [WIDTH - 1 : 0] operand_1,
    input wire [WIDTH - 1 : 0] operand_2,
    
    input wire [ 1 : 0] operation,

    output reg [WIDTH - 1 : 0] result,
    output reg ready
);

    always @(*)
    begin
        case (operation)
            `FPU_ADD    : begin result <= operand_1 + operand_2; ready <= 1; end
            `FPU_SUB    : begin result <= operand_1 - operand_2; ready <= 1; end
            `FPU_MUL    : begin result <= product[WIDTH + FBITS - 1 : FBITS]; ready <= product_ready; end
            `FPU_SQRT   : begin result <= root; ready <= root_ready; end
            default     : begin result <= 'bz; ready <= 0; end
        endcase
    end

    always @(posedge reset)
    begin
        if (reset)  ready = 0;
        else        ready = 'bz;
    end
    // ------------------- //
    // Square Root Circuit //
    // ------------------- //
    reg [WIDTH - 1 : 0] root;
    reg root_ready;

    reg [3:0] sqrt_state;
    reg [WIDTH - 1 : 0] radicand;
    reg [WIDTH - 1 : 0] res;
    reg [WIDTH - 1 : 0] iteration;
    reg [WIDTH - 1 : 0] temp;
    reg [WIDTH - 1 : 0] reminder;
    reg [WIDTH - 1 : 0] op1;
    reg [1 : 0] bits;

    always @(posedge clk or posedge reset)
    begin
        if (reset) begin
            sqrt_state <=0;
            root <= 0;
            root_ready <= 0;
            op1 <= operand_1;
        end else if (operation == `FPU_SQRT) begin
            case (sqrt_state)
                0: begin // Initialize
                    radicand <= operand_1[WIDTH - 1: WIDTH - 2];
                    res <= 0;
                    temp <= 2'b01;
                    sqrt_state <= 1;
                    iteration <= (WIDTH + FBITS) / 2;
                end
                1: begin // Main calculation loop
                    if(iteration > 0) begin
                        reminder <= radicand - temp;
                        if(reminder < 0) begin
                            res = res << 1;
                        end else begin
                            res = (res << 1) + 1;
                        end
                    end
                    
                    op1 <= op1 << 2;
                    bits <= op1[WIDTH - 1 : WIDTH - 2];
                    radicand <= (radicand << 2) + bits;
                    temp <= (res << 2) + 1 ;    
                    iteration <= iteration - 1;

                end
                2: begin // Set ready signal
                    root <= res;
                    root_ready <= 1;
                    sqrt_state <= 0;
                end
            endcase
        end    
    end

    
        /*
         *  Describe Your Square Root Calculator Circuit Here.
         */

    // ------------------ //
    // Multiplier Circuit //
    // ------------------ //   
    reg [64 - 1 : 0] product;
    reg product_ready;

    reg     [15 : 0] multiplierCircuitInput1;
    reg     [15 : 0] multiplierCircuitInput2;
    wire    [31 : 0] multiplierCircuitResult;

    Multiplier multiplier_circuit
    (
        .operand_1(multiplierCircuitInput1),
        .operand_2(multiplierCircuitInput2),
        .product(multiplierCircuitResult)
    );

    reg     [31 : 0] partialProduct1;
    reg     [31 : 0] partialProduct2;
    reg     [31 : 0] partialProduct3;
    reg     [31 : 0] partialProduct4;
    
    reg[2:0] mul_state;

    always @(posedge clk or posedge reset)
    begin
        if (reset) begin
            product <= 0;
            mul_state <= 0;
            product_ready <= 0;
        end else if (operation == `FPU_MUL) begin
            case (mul_state)
                0: begin // Start LL multiplication
                    multiplierCircuitInput1 <= operand_1[15:0];
                    multiplierCircuitInput2 <= operand_2[15:0];
                    mul_state <= 1;
                end
                1: begin // LL multiplication done, start LH
                    partialProduct1 <= multiplierCircuitResult;
                    multiplierCircuitInput1 <= operand_1[15:0];
                    multiplierCircuitInput2 <= operand_2[31:16];
                    mul_state <= 2;
                end
                2: begin // LH multiplication done, start HL
                    partialProduct2 <= multiplierCircuitResult << 16;
                    multiplierCircuitInput1 <= operand_1[31:16];
                    multiplierCircuitInput2 <= operand_2[15:0];
                    mul_state <= 3;
                end
                3: begin // HL multiplication done, start HH
                    partialProduct3 <= multiplierCircuitResult << 16;
                    multiplierCircuitInput1 <= operand_1[31:16];
                    multiplierCircuitInput2 <= operand_2[31:16];
                    mul_state <= 4;
                end
                4: begin // HH multiplication done, combine results
                    partialProduct4 <= multiplierCircuitResult << 32;
                    mul_state <= 5;
                end
                5: begin 
                    product <= partialProduct4 + partialProduct3 + partialProduct2 + partialProduct1;
                    product_ready <= 1;
                end
                default: mul_state <= 0;
            endcase
        end
    end
        /*
         *  Describe Your 32-bit Multiplier Circuit Here.
         */
         
endmodule

module Multiplier
(
    input wire [15 : 0] operand_1,
    input wire [15 : 0] operand_2,

    output reg [31 : 0] product
);

    always @(*)
    begin
        product <= operand_1 * operand_2;
    end
endmodule